-------------------------------------------------------------------------------
-- Design: FSM LED Shifting                                                  --
--                                                                           --
-- Author : Sebastian Dichler                                                --
-- Date : 15 Oktober 2017                                                    --
-- File : tb_fsm_led_shift.vhd                                                        --
-------------------------------------------------------------------------------

